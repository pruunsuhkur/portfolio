module lut_based_nco #( parameter LUT_WIDTH  = 16, 
                                  LUT_LENGTH = 6, 
                       localparam PHASE_BITWIDTH_INTEGER = LUT_LENGTH, 
                                  PHASE_BITWIDTH_FRACTIONAL = 2, 
                                  ACC_SIZE = PHASE_BITWIDTH_INTEGER + PHASE_BITWIDTH_FRACTIONAL)
(
    input  wire                              iclk, 
    input  wire                              iresetn,
    input  wire       [ACC_SIZE + 1 - 1 : 0] step,
    output reg signed [LUT_WIDTH    - 1 : 0] out 
);
    
    reg [ACC_SIZE   + 1 : 0] accum; 
    reg [LUT_WIDTH  - 1 : 0] LUT [2**LUT_LENGTH - 1 : 0]; 
    
    always @(posedge iclk or negedge iresetn)
        if (~iresetn)
            begin
                LUT[ 0] <= 16'b000000000000000; 
                LUT[ 1] <= 16'b000000000000000; 
                LUT[ 2] <= 16'b000000000000000; 
                LUT[ 3] <= 16'b000000000000000; 
                LUT[ 4] <= 16'b000000000000000; 
                LUT[ 5] <= 16'b000000000000000; 
                LUT[ 6] <= 16'b000000000000000; 
                LUT[ 7] <= 16'b000000000000000; 
                LUT[ 8] <= 16'b000000000000000; 
                LUT[ 9] <= 16'b000000000000000; 
                LUT[10] <= 16'b000000000000000; 
                LUT[11] <= 16'b000000000000000; 
                LUT[12] <= 16'b000000000000000; 
                LUT[13] <= 16'b000000000000000; 
                LUT[14] <= 16'b000000000000000; 
                LUT[15] <= 16'b000000000000000; 
                LUT[16] <= 16'b000000000000000; 
                LUT[17] <= 16'b000000000000000; 
                LUT[18] <= 16'b000000000000000; 
                LUT[19] <= 16'b000000000000000; 
                LUT[20] <= 16'b000000000000000; 
                LUT[21] <= 16'b000000000000000; 
                LUT[22] <= 16'b000000000000000; 
                LUT[23] <= 16'b000000000000000; 
                LUT[24] <= 16'b000000000000000; 
                LUT[25] <= 16'b000000000000000; 
                LUT[26] <= 16'b000000000000000; 
                LUT[27] <= 16'b000000000000000; 
                LUT[28] <= 16'b000000000000000; 
                LUT[29] <= 16'b000000000000000; 
                LUT[30] <= 16'b000000000000000; 
                LUT[31] <= 16'b000000000000000; 
                LUT[32] <= 16'b000000000000000; 
                LUT[33] <= 16'b000000000000000; 
                LUT[34] <= 16'b000000000000000; 
                LUT[35] <= 16'b000000000000000; 
                LUT[36] <= 16'b000000000000000; 
                LUT[37] <= 16'b000000000000000; 
                LUT[38] <= 16'b000000000000000; 
                LUT[39] <= 16'b000000000000000; 
                LUT[40] <= 16'b000000000000000; 
                LUT[41] <= 16'b000000000000000; 
                LUT[42] <= 16'b000000000000000; 
                LUT[43] <= 16'b000000000000000; 
                LUT[44] <= 16'b000000000000000; 
                LUT[45] <= 16'b000000000000000; 
                LUT[46] <= 16'b000000000000000; 
                LUT[47] <= 16'b000000000000000; 
                LUT[48] <= 16'b000000000000000; 
                LUT[49] <= 16'b000000000000000; 
                LUT[50] <= 16'b000000000000000; 
                LUT[51] <= 16'b000000000000000; 
                LUT[52] <= 16'b000000000000000; 
                LUT[53] <= 16'b000000000000000; 
                LUT[54] <= 16'b000000000000000; 
                LUT[55] <= 16'b000000000000000; 
                LUT[56] <= 16'b000000000000000; 
                LUT[57] <= 16'b000000000000000; 
                LUT[58] <= 16'b000000000000000; 
                LUT[59] <= 16'b000000000000000; 
                LUT[60] <= 16'b000000000000000; 
                LUT[61] <= 16'b000000000000000; 
                LUT[62] <= 16'b000000000000000; 
                LUT[63] <= 16'b000000000000000; 
            end
        else
            begin
                LUT[ 0] <= 16'b0000000000000000; 
                LUT[ 1] <= 16'b0000001100101010; 
                LUT[ 2] <= 16'b0000011001010100; 
                LUT[ 3] <= 16'b0000100101111101; 
                LUT[ 4] <= 16'b0000110010100101; 
                LUT[ 5] <= 16'b0000111111001010; 
                LUT[ 6] <= 16'b0001001011101101; 
                LUT[ 7] <= 16'b0001011000001101; 
                LUT[ 8] <= 16'b0001100100101010; 
                LUT[ 9] <= 16'b0001110001000011; 
                LUT[10] <= 16'b0001111101010111; 
                LUT[11] <= 16'b0010001001100110; 
                LUT[12] <= 16'b0010010101110000; 
                LUT[13] <= 16'b0010100001110100; 
                LUT[14] <= 16'b0010101101110010; 
                LUT[15] <= 16'b0010111001101001; 
                LUT[16] <= 16'b0011000101011001; 
                LUT[17] <= 16'b0011010001000001; 
                LUT[18] <= 16'b0011011100100001; 
                LUT[19] <= 16'b0011100111111000; 
                LUT[20] <= 16'b0011110011000110; 
                LUT[21] <= 16'b0011111110001010; 
                LUT[22] <= 16'b0100001001000101; 
                LUT[23] <= 16'b0100010011110101; 
                LUT[24] <= 16'b0100011110011011; 
                LUT[25] <= 16'b0100101000110101; 
                LUT[26] <= 16'b0100110011000011; 
                LUT[27] <= 16'b0100111101000110; 
                LUT[28] <= 16'b0101000110111100; 
                LUT[29] <= 16'b0101010000100101; 
                LUT[30] <= 16'b0101011010000010; 
                LUT[31] <= 16'b0101100011010000; 
                LUT[32] <= 16'b0101101100010001; 
                LUT[33] <= 16'b0101110101000011; 
                LUT[34] <= 16'b0101111101100111; 
                LUT[35] <= 16'b0110000101111100; 
                LUT[36] <= 16'b0110001110000010; 
                LUT[37] <= 16'b0110010101111000; 
                LUT[38] <= 16'b0110011101011110; 
                LUT[39] <= 16'b0110100100110100; 
                LUT[40] <= 16'b0110101011111001; 
                LUT[41] <= 16'b0110110010101110; 
                LUT[42] <= 16'b0110111001010001; 
                LUT[43] <= 16'b0110111111100100; 
                LUT[44] <= 16'b0111000101100101; 
                LUT[45] <= 16'b0111001011010100; 
                LUT[46] <= 16'b0111010000110001; 
                LUT[47] <= 16'b0111010101111100; 
                LUT[48] <= 16'b0111011010110100; 
                LUT[49] <= 16'b0111011111011010; 
                LUT[50] <= 16'b0111100011101101; 
                LUT[51] <= 16'b0111100111101101; 
                LUT[52] <= 16'b0111101011011011; 
                LUT[53] <= 16'b0111101110110100; 
                LUT[54] <= 16'b0111110001111011; 
                LUT[55] <= 16'b0111110100101110; 
                LUT[56] <= 16'b0111110111001101; 
                LUT[57] <= 16'b0111111001011001; 
                LUT[58] <= 16'b0111111011010001; 
                LUT[59] <= 16'b0111111100110101; 
                LUT[60] <= 16'b0111111110000101; 
                LUT[61] <= 16'b0111111111000001; 
                LUT[62] <= 16'b0111111111101001; 
                LUT[63] <= 16'b0111111111111101; 
            end
    
    always @(posedge iclk or negedge iresetn) 
        if (~iresetn)
            accum <= 10'b0;
        else 
            accum <= accum  + step;
          
    always @(posedge iclk or negedge iresetn) 
        if (~iresetn)
            out <= 16'b0;
        else
            case (accum[ACC_SIZE + 1 : ACC_SIZE])
                2'b00: out <=  LUT[ accum[ACC_SIZE - 1 : PHASE_BITWIDTH_FRACTIONAL]];
                2'b01: out <=  LUT[~accum[ACC_SIZE - 1 : PHASE_BITWIDTH_FRACTIONAL]];
                2'b10: out <= ~LUT[ accum[ACC_SIZE - 1 : PHASE_BITWIDTH_FRACTIONAL]];
                2'b11: out <= ~LUT[~accum[ACC_SIZE - 1 : PHASE_BITWIDTH_FRACTIONAL]];
            endcase

endmodule
